** Profile: "SCHEMATIC1-sim1"  [ C:\Users\Justin\Documents\School\2024-2025\Fall Quarter\EEC 100\OrCAD Lab Simulations\EEC-100-OrCAD-Simulations\lab 8-laplace transform analysis-PSpiceFiles\SCHEMATIC1\sim1.sim ] 

** Creating circuit file "sim1.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Profile Libraries :
* Local Libraries :
* From [PSPICE NETLIST] section of C:\Users\Justin\AppData\Roaming\SPB_Data\cdssetup\OrCAD_PSpice\17.2.0\PSpice.ini file:
.lib "nomd.lib" 

*Analysis directives: 
.TRAN  0 6ms 0 1u 
.OPTIONS ADVCONV
.PROBE64 V(alias(*)) I(alias(*)) W(alias(*)) D(alias(*)) NOISE(alias(*)) 
.INC "..\SCHEMATIC1.net" 


.END
